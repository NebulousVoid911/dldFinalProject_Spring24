module game(input clk, reset, d, seed, shift_seed, d0, d1, s,   output q, y);

flopr flopr1();



mux2 select();



lfsr64 randomizer();



endmodule