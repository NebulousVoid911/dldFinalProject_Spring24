module game(input clk, reset, d, seed, shift_seed,  output q);

flopr flopr1();



mux2 select();



lfsr64 randomizer();



endmodule